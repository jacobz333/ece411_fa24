module plru_logic (
    
);

endmodule