/*
 * decodes the given instruction 
 * 
 */
module decode_logic #(
    parameter   PR_BITS       = 5,
    localparam  PR_NUM        = 2**PR_BITS,
    parameter   ROBSIZE_BITS  = 4
) (

);

endmodule
